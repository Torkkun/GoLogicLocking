module test_module (A, B, C, D);
//no parameter
  input A
  input B
  input C
  output D
//no register decl
//no event decl
//no net decl
//no premitive decl
endmodule